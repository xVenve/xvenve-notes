* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\Sesion0\C7.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 29 16:46:40 2019



** Analysis setup **
.tran 0 2
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "C7.net"
.INC "C7.als"


.probe


.END
