* F:\PSPICE\Sesion0\C1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 17 13:01:11 2019



** Analysis setup **
.DC LIN V_V1 0 200 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "C1.net"
.INC "C1.als"


.probe


.END
