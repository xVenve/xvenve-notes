* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\Sesion0\C3.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 29 15:41:26 2019



** Analysis setup **
.DC LIN  0 20 1 
.tran 0ns 1000ns SKIPBP
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "C3.net"
.INC "C3.als"


.probe


.END
