* F:\PSPICE\Sesion0\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 17 12:46:22 2019



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
