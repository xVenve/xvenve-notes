* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\P1\Ej1.2.sch

* Schematics Version 9.1 - Web Update 1
* Mon Apr 08 17:55:24 2019



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ej1.2.net"
.INC "Ej1.2.als"


.probe


.END
