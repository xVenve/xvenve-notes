* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\P1\Ej3.2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Apr 12 18:44:21 2019



** Analysis setup **
.DC LIN V_V3 0 400 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ej3.2.net"
.INC "Ej3.2.als"


.probe


.END
