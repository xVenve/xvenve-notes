* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\Sesion0\C6.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 29 16:33:12 2019



** Analysis setup **
.tran 0ns 10 SKIPBP
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "C6.net"
.INC "C6.als"


.probe


.END
