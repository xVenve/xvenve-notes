* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\Sesion0\C4.sch

* Schematics Version 9.1 - Web Update 1
* Fri Mar 29 16:10:22 2019



** Analysis setup **
.tran 0 20 SKIPBP
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "C4.net"
.INC "C4.als"


.probe


.END
