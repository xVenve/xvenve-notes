* W:\Universidad\Primero\2�. Cuatrimestre\PRINCIPIOS FISICOS DE LA INGENIER�A INFORMATICA\PSPICE\P1\Ej6.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 11 19:11:02 2019



** Analysis setup **
.tran 0 8ms SKIPBP
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ej6.net"
.INC "Ej6.als"


.probe


.END
